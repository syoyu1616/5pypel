`include "define.v"

module writeback(
    input rst,
    input clk,
    input keep, //nopとかのときに一緒に使うやつでpcの維持など
    input nop,

    input [31:0] PCp4_pype3,
    input [31:0] mem_data_pype,
    input [31:0] ALU_co_pype3,
    input [4:0] WReg_pype3,

    input RegWrite_pype3,
    input [1:0]MemtoReg_pype3,

    input [1:0] ID_EX_write_pype3,
    input [1:0] ID_EX_write_addi_pype3,
    input [1:0] forwarding_stall_load_pyc_pype3,


    output  [31:0] write_reg_data,
    output  Regwrite,
    output  [4:0] write_reg_address,
    output  [1:0] ID_EX_write,
    output  [1:0] ID_EX_write_addi,
    output  [1:0] forwarding_stall_load_pyc
);

assign write_reg_data = 
        MemtoReg_pype3 == `write_reg_PCp4 ? PCp4_pype3 : //jalrのシングルラインの場合　パイプラインの場合mucを012まで増やすことを考慮
        MemtoReg_pype3 == `write_reg_memd ? mem_data_pype : ALU_co_pype3;

assign Regwrite = ~RegWrite_pype3;

assign write_reg_address = WReg_pype3;

assign ID_EX_write = ID_EX_write_pype3;
assign ID_EX_write_addi = ID_EX_write_addi_pype3;
assign forwarding_stall_load_pyc = forwarding_stall_load_pyc_pype3;
//memtoregの伝達が途中で止まってるせいでwriteが上手くいってない


endmodule